`ifndef STAGE1_CONTROL
`define STAGE1_CONTROL

// PC_Mux Control
`define PC_SEL_PC_4      1'b0
`define PC_SEL_ALU_OUT   1'b1

`endif //STAGE1_CONTROL