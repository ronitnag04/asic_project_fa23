`ifndef MWControl
`define MWControl

// wb_sel
`define SEL_MEM         2'd0
`define SEL_ALU         2'd1
`define SEL_PC4         2'd2

`endif //MWControl